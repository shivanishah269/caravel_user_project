VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN L1_hit_count[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END L1_hit_count[0]
  PIN L1_hit_count[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.920 900.000 300.520 ;
    END
  END L1_hit_count[1]
  PIN L1_hit_count[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END L1_hit_count[2]
  PIN L1_hit_count[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 596.000 150.330 600.000 ;
    END
  END L1_hit_count[3]
  PIN L1_hit_count[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 596.000 450.250 600.000 ;
    END
  END L1_hit_count[4]
  PIN L1_hit_count[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END L1_hit_count[5]
  PIN L1_hit_count[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END L1_hit_count[6]
  PIN L1_hit_count[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END L1_hit_count[7]
  PIN L1_hit_count[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END L1_hit_count[8]
  PIN L1_hit_count[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 596.000 750.170 600.000 ;
    END
  END L1_hit_count[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 6.990 595.720 149.770 596.090 ;
        RECT 150.610 595.720 449.690 596.090 ;
        RECT 450.530 595.720 749.610 596.090 ;
        RECT 750.450 595.720 890.470 596.090 ;
        RECT 6.990 4.280 890.470 595.720 ;
        RECT 6.990 4.000 74.790 4.280 ;
        RECT 75.630 4.000 224.750 4.280 ;
        RECT 225.590 4.000 374.710 4.280 ;
        RECT 375.550 4.000 524.670 4.280 ;
        RECT 525.510 4.000 674.630 4.280 ;
        RECT 675.470 4.000 824.590 4.280 ;
        RECT 825.430 4.000 890.470 4.280 ;
      LAYER met3 ;
        RECT 4.000 450.520 896.000 587.685 ;
        RECT 4.400 449.120 896.000 450.520 ;
        RECT 4.000 300.920 896.000 449.120 ;
        RECT 4.000 299.520 895.600 300.920 ;
        RECT 4.000 150.640 896.000 299.520 ;
        RECT 4.400 149.240 896.000 150.640 ;
        RECT 4.000 10.715 896.000 149.240 ;
      LAYER met4 ;
        RECT 334.255 222.535 404.640 422.785 ;
        RECT 407.040 222.535 481.440 422.785 ;
        RECT 483.840 222.535 558.240 422.785 ;
        RECT 560.640 222.535 562.745 422.785 ;
  END
END user_proj_example
END LIBRARY


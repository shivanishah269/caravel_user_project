magic
tech sky130A
magscale 1 2
timestamp 1641881671
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 30010 119200 30066 120000
rect 89994 119200 90050 120000
rect 149978 119200 150034 120000
rect 15014 0 15070 800
rect 45006 0 45062 800
rect 74998 0 75054 800
rect 104990 0 105046 800
rect 134982 0 135038 800
rect 164974 0 165030 800
<< obsm2 >>
rect 1398 119144 29954 119218
rect 30122 119144 89938 119218
rect 90106 119144 149922 119218
rect 150090 119144 178094 119218
rect 1398 856 178094 119144
rect 1398 800 14958 856
rect 15126 800 44950 856
rect 45118 800 74942 856
rect 75110 800 104934 856
rect 105102 800 134926 856
rect 135094 800 164918 856
rect 165086 800 178094 856
<< metal3 >>
rect 0 89904 800 90024
rect 179200 59984 180000 60104
rect 0 29928 800 30048
<< obsm3 >>
rect 800 90104 179200 117537
rect 880 89824 179200 90104
rect 800 60184 179200 89824
rect 800 59904 179120 60184
rect 800 30128 179200 59904
rect 880 29848 179200 30128
rect 800 2143 179200 29848
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 66851 44507 80928 84557
rect 81408 44507 96288 84557
rect 96768 44507 111648 84557
rect 112128 44507 112549 84557
<< labels >>
rlabel metal3 s 0 89904 800 90024 6 L1_hit_count[0]
port 1 nsew signal output
rlabel metal3 s 179200 59984 180000 60104 6 L1_hit_count[1]
port 2 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 L1_hit_count[2]
port 3 nsew signal output
rlabel metal2 s 30010 119200 30066 120000 6 L1_hit_count[3]
port 4 nsew signal output
rlabel metal2 s 89994 119200 90050 120000 6 L1_hit_count[4]
port 5 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 L1_hit_count[5]
port 6 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 L1_hit_count[6]
port 7 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 L1_hit_count[7]
port 8 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 L1_hit_count[8]
port 9 nsew signal output
rlabel metal2 s 149978 119200 150034 120000 6 L1_hit_count[9]
port 10 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 clk
port 11 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 reset
port 12 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 14 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 15460442
string GDS_START 427542
<< end >>

